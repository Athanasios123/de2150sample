LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY comparator IS
PORT ( 
   C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	Z : OUT STD_LOGIC
	);
END comparator;

ARCHITECTURE comparator_arch OF comparator IS
BEGIN
process(C)
	begin
		case C is
			when "0000" =>   Z <= '0';-- 0
			when "0001" =>   Z <= '0';-- 0
			when "0010" =>   Z <= '0';-- 0
			when "0011" =>   Z <= '0';-- 0
			when "0100" =>   Z <= '0';-- 0
			when "0101" =>   Z <= '0';-- 0
			when "0110" =>   Z <= '0';-- 0
			when "0111" =>   Z <= '0';-- 0
			when "1000" =>   Z <= '0';-- 0
			when "1001" =>   Z <= '0';-- 0
         when others => Z <= '1';-- 
		end case;
end process;
END comparator_arch;